two_stage_amp power supply gain test

* Two stage OPAMP
.include "{{include}}"
.param wp1=0.5u lp1=90n mp1={{mp1}}
.param wn1=0.5u ln1=90n mn1={{mn1}}
.param wn3=0.5u ln3=90n mn3={{mn3}}
.param wp3=0.5u lp3=90n mp3={{mp3}}
.param wn4=0.5u ln4=90n mn4={{mn4}}
.param wn5=0.5u ln5=90n mn5={{mn5}}
.param cc={{cc}}
.param rz={{rz}}
.param ibias=30u
.param cload=10p
.param vcm=0.6

* parasitic modeling
cpar_out net6 VSS {(mn5+mp3) * 5f + rz * 1f}
cpar8 net8 VSS {cc * 0.05 + rz * 1f}
cpar_o1 net5 VSS {cc * 0.03 + (mp1 + mn1 + mp3) * 5f}
cpar_m net4 VSS {(2 * mp1 + mn1) * 5f}
cpar_tail net3 VSS {(2 * mn1 + mn3) * 5f}
cpar_bias net7 VSS {(mn4 + mn3 + mn5) * 5f}

mp1 net4 net4 VDD VDD pmos w=wp1 l=lp1 m=mp1
mp2 net5 net4 VDD VDD pmos w=wp1 l=lp1 m=mp1
mn1 net4 net2 net3 net3 nmos w=wn1 l=ln1 m=mn1
mn2 net5 net1 net3 net3 nmos w=wn1 l=ln1 m=mn1
mn3 net3 net7 VSS VSS nmos w=wn3 l=ln3 m=mn3
mn4 net7 net7 VSS VSS nmos w=wn4 l=ln4 m=mn4
mp3 net6 net5 VDD VDD pmos w=wp3 l=lp3 m=mp3
mn5 net6 net7 VSS VSS nmos w=wn5 l=ln5 m=mn5
cc net5 net8 cc
rz net8 net6 rz
ibias VDD net7 ibias

vin in 0 dc=0 ac=0
ein1 net1 cm in 0 0.5
ein2 net2 cm in 0 -0.5
vcm cm 0 dc=vcm

vindd VDD_dc VDD ac=1
vdd VDD_dc 0 dc=1.2
vss 0 VSS dc=0
CL net6 0 cload

.ac dec 10 1 10G

.control
run
set units=degrees
set wr_vecnames
option numdgt=7
wrdata {{ps}} v(net6)
.endc

.end
